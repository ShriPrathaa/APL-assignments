.circuit
V1   2 1  dc 20
V2   4   3  dc   10
I1    GND 2  dc   10
R1 1 4 1
R2 2 3 2
R3 4 GND 3
R4 1 GND 4
R5 3 GND 5
.end