.circuit
V1   1 GND  dc 2
R1   1   2     1
R2   2 GND     1
V3 1 5 dc 6
.end