.circuit
V3 GND 1 dc 10
V1 GND 2 dc 5
V2 GND 3 dc 2
R1 2 3 2
R2  1 3  1
R3  1 2  3
.end